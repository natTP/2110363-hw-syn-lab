`timescale 1ns / 1ps
//-------------------------------------------------------
// File name    : nano_sc_system.v
// Title        : nanoCPU Single Cycle system.
// Library      : nanoLADA
// Purpose      : Computer Architecture
// Developers   : Krerk Piromsopa, Ph. D.
//              : Chulalongkorn University.

module nano_sc_system(
);
wire 	[31:0]	p_address;
wire 	[31:0]	p_data;
wire	[31:0]	d_address;
wire		mem_wr;
wire	[31:0]	d_data;
reg		clk;
reg		nreset;

nanocpu	CPU(p_address,p_data,d_address,d_data,mem_wr,clk,nreset);
rom 	PROGMEM(p_data,p_address[17:2]);
memory 	DATAMEM(d_data,d_address[15:0],mem_wr,clk,sw,seg,an,dp);

initial
begin
	$dumpfile("nano_sc_system.dump");
	$dumpvars(4, nano_sc_system);

	clk=0;
	nreset=0;
	#100;
	nreset=1;
	#2000;
	$finish;
end

always
begin : CLOCK
	#20
	clk=~clk;
end


endmodule
